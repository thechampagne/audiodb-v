/*
 * Copyright 2022 XXIV
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */
module model

pub struct Artist {
pub:
	id_artist           string [json: idArtist]
	str_artist          string [json: strArtist]
	str_artiststripped  string [json: strArtistStripped]
	str_artistalternate string [json: strArtistAlternate]
	str_label           string [json: strLabel]
	id_label            string [json: idLabel]
	int_formedyear      string [json: intFormedYear]
	int_bornyear        string [json: intBornYear]
	int_diedyear        string [json: intDiedYear]
	str_disbanded       string [json: strDisbanded]
	str_style           string [json: strStyle]
	str_genre           string [json: strGenre]
	str_mood            string [json: strMood]
	str_website         string [json: strWebsite]
	str_facebook        string [json: strFacebook]
	str_twitter         string [json: strTwitter]
	str_biographyen     string [json: strBiographyEN]
	str_biographyde     string [json: strBiographyDE]
	str_biographyfr     string [json: strBiographyFR]
	str_biographycn     string [json: strBiographyCN]
	str_biographyit     string [json: strBiographyIT]
	str_biographyjp     string [json: strBiographyJP]
	str_biographyru     string [json: strBiographyRU]
	str_biographyes     string [json: strBiographyES]
	str_biographypt     string [json: strBiographyPT]
	str_biographyse     string [json: strBiographySE]
	str_biographynl     string [json: strBiographyNL]
	str_biographyhu     string [json: strBiographyHU]
	str_biographyno     string [json: strBiographyNO]
	str_biographyil     string [json: strBiographyIL]
	str_biographypl     string [json: strBiographyPL]
	str_gender          string [json: strGender]
	int_members         string [json: intMembers]
	str_country         string [json: strCountry]
	str_countrycode     string [json: strCountryCode]
	str_artistthumb     string [json: strArtistThumb]
	str_artistlogo      string [json: strArtistLogo]
	str_artistcutout    string [json: strArtistCutout]
	str_artistclearart  string [json: strArtistClearart]
	str_artistwidethumb string [json: strArtistWideThumb]
	str_artistfanart    string [json: strArtistFanart]
	str_artistfanart2   string [json: strArtistFanart2]
	str_artistfanart3   string [json: strArtistFanart3]
	str_artistfanart4   string [json: strArtistFanart4]
	str_artistbanner    string [json: strArtistBanner]
	str_musicbrainzid   string [json: strMusicBrainzID]
	str_isnicode        string [json: strISNIcode]
	str_lastfmchart     string [json: strLastFMChart]
	int_charted         string [json: intCharted]
	str_locked          string [json: strLocked]
}

pub struct Discography {
pub:
	str_album         string [json: strAlbum]
	int_year_released string [json: intYearReleased]
}

pub struct Album {
pub:
	id_album                string [json: idAlbum]
	id_artist               string [json: idArtist]
	id_label                string [json: idLabel]
	str_album               string [json: strAlbum]
	str_albumstripped       string [json: strAlbumStripped]
	str_artist              string [json: strArtist]
	str_artiststripped      string [json: strArtistStripped]
	int_yearreleased        string [json: intYearReleased]
	str_style               string [json: strStyle]
	str_genre               string [json: strGenre]
	str_label               string [json: strLabel]
	str_releaseformat       string [json: strReleaseFormat]
	int_sales               string [json: intSales]
	str_albumthumb          string [json: strAlbumThumb]
	str_albumthumbhq        string [json: strAlbumThumbHQ]
	str_albumthumbback      string [json: strAlbumThumbBack]
	str_albumcdart          string [json: strAlbumCDart]
	str_albumspine          string [json: strAlbumSpine]
	str_album3dcase         string [json: strAlbum3DCase]
	str_album3dflat         string [json: strAlbum3DFlat]
	str_album3dface         string [json: strAlbum3DFace]
	str_album3dthumb        string [json: strAlbum3DThumb]
	str_descriptionen       string [json: strDescriptionEN]
	str_descriptionde       string [json: strDescriptionDE]
	str_descriptionfr       string [json: strDescriptionFR]
	str_descriptioncn       string [json: strDescriptionCN]
	str_descriptionit       string [json: strDescriptionIT]
	str_descriptionjp       string [json: strDescriptionJP]
	str_descriptionru       string [json: strDescriptionRU]
	str_descriptiones       string [json: strDescriptionES]
	str_descriptionpt       string [json: strDescriptionPT]
	str_descriptionse       string [json: strDescriptionSE]
	str_descriptionnl       string [json: strDescriptionNL]
	str_descriptionhu       string [json: strDescriptionHU]
	str_descriptionno       string [json: strDescriptionNO]
	str_descriptionil       string [json: strDescriptionIL]
	str_descriptionpl       string [json: strDescriptionPL]
	int_loved               string [json: intLoved]
	int_score               string [json: intScore]
	int_scorevotes          string [json: intScoreVotes]
	str_review              string [json: strReview]
	str_mood                string [json: strMood]
	str_theme               string [json: strTheme]
	str_speed               string [json: strSpeed]
	str_location            string [json: strLocation]
	str_musicbrainzid       string [json: strMusicBrainzID]
	str_musicbrainzartistid string [json: strMusicBrainzArtistID]
	str_allmusicid          string [json: strAllMusicID]
	str_bbcreviewid         string [json: strBBCReviewID]
	str_rateyourmusicid     string [json: strRateYourMusicID]
	str_discogsid           string [json: strDiscogsID]
	str_wikidataid          string [json: strWikidataID]
	str_wikipediaid         string [json: strWikipediaID]
	str_geniusid            string [json: strGeniusID]
	str_lyricwikiid         string [json: strLyricWikiID]
	str_musicmozid          string [json: strMusicMozID]
	str_itunesid            string [json: strItunesID]
	str_amazonid            string [json: strAmazonID]
	str_locked              string [json: strLocked]
}

pub struct Track {
pub:
	id_track                string [json: idTrack]
	id_album                string [json: idAlbum]
	id_artist               string [json: idArtist]
	id_lyric                string [json: idLyric]
	id_imvdb                string [json: idIMVDB]
	str_track               string [json: strTrack]
	str_album               string [json: strAlbum]
	str_artist              string [json: strArtist]
	str_artistalternate     string [json: strArtistAlternate]
	int_cd                  string [json: intCD]
	int_duration            string [json: intDuration]
	str_genre               string [json: strGenre]
	str_mood                string [json: strMood]
	str_style               string [json: strStyle]
	str_theme               string [json: strTheme]
	str_descriptionen       string [json: strDescriptionEN]
	str_descriptionde       string [json: strDescriptionDE]
	str_descriptionfr       string [json: strDescriptionFR]
	str_descriptioncn       string [json: strDescriptionCN]
	str_descriptionit       string [json: strDescriptionIT]
	str_descriptionjp       string [json: strDescriptionJP]
	str_descriptionru       string [json: strDescriptionRU]
	str_descriptiones       string [json: strDescriptionES]
	str_descriptionpt       string [json: strDescriptionPT]
	str_descriptionse       string [json: strDescriptionSE]
	str_descriptionnl       string [json: strDescriptionNL]
	str_descriptionhu       string [json: strDescriptionHU]
	str_descriptionno       string [json: strDescriptionNO]
	str_descriptionil       string [json: strDescriptionIL]
	str_descriptionpl       string [json: strDescriptionPL]
	str_trackthumb          string [json: strTrackThumb]
	str_track3dcase         string [json: strTrack3DCase]
	str_tracklyrics         string [json: strTrackLyrics]
	str_musicvid            string [json: strMusicVid]
	str_musicviddirector    string [json: strMusicVidDirector]
	str_musicvidcompany     string [json: strMusicVidCompany]
	str_musicvidscreen1     string [json: strMusicVidScreen1]
	str_musicvidscreen2     string [json: strMusicVidScreen2]
	str_musicvidscreen3     string [json: strMusicVidScreen3]
	int_musicvidviews       string [json: intMusicVidViews]
	int_musicvidlikes       string [json: intMusicVidLikes]
	int_musicviddislikes    string [json: intMusicVidDislikes]
	int_musicvidfavorites   string [json: intMusicVidFavorites]
	int_musicvidcomments    string [json: intMusicVidComments]
	int_tracknumber         string [json: intTrackNumber]
	int_loved               string [json: intLoved]
	int_score               string [json: intScore]
	int_scorevotes          string [json: intScoreVotes]
	int_totallisteners      string [json: intTotalListeners]
	int_totalplays          string [json: intTotalPlays]
	str_musicbrainzid       string [json: strMusicBrainzID]
	str_musicbrainzalbumid  string [json: strMusicBrainzAlbumID]
	str_musicbrainzartistid string [json: strMusicBrainzArtistID]
	str_locked              string [json: strLocked]
}

pub struct MusicVideo {
pub:
	id_artist         string [json: idArtist]
	id_album          string [json: idAlbum]
	id_track          string [json: idTrack]
	str_track         string [json: strTrack]
	str_trackthumb    string [json: strTrackThumb]
	str_musicvid      string [json: strMusicVid]
	str_descriptionen string [json: strDescriptionEN]
}
